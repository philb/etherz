module data_fifo();
   reg [7:0] data;
   reg [7:0] data_next;   

   reg 	     data_full;
   reg 	     data_next_full;   
   
endmodule // data_fifo
