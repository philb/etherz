module taskfile();
   
   reg [7:0] command;
   reg [7:0] lba0;
   reg [7:0] lba1;
   reg [7:0] lba2;
   reg [7:0] lba3;
   reg [7:0] sector_count;   
   reg [7:0] status;

endmodule // taskfile
